library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;
use IEEE.std_logic_textio.all;
use std.env.all;

use work.param_disenyo_pkg.all;
use work.camino_dat_pkg.all;
use work.peticiones_cache_pkg.all;
use work.controlador_pkg.all;

use work.procedimientos_peticiones_pkg.all;

use work.impri_memoria_pkg.all;
use work.impri_cache_pkg.all;
--use work.impri_traza_pkg.all;

entity prueba_ensamblado is
    generic(pasoapaso: integer range 0 to 1:= 0;
			   imprimir_traza: integer:= 0;
			   imprimir_CACHE: integer:= 1;
			   imprimir_MEMORIA: integer:= 1;
			   comprobar_load: integer:= 1);
end prueba_ensamblado;
  
architecture prueba of prueba_ensamblado is

component jerarquia is 
 port(reloj: in std_logic;
      pcero: in std_logic;
		pet_proc: in tp_peticion; 
		resp_cache: out tp_respuesta;
		cache_lista: out std_logic);
end component;

signal reloj, pcero: std_logic;

signal peticion: tp_peticion;
signal respuesta: tp_respuesta;
signal pet_listo: std_logic;

signal s_mem_etiq: tp_m_ET;
signal s_mem_estado: tp_m_EST;
signal s_mem_datos: tp_m_DAT;
signal s_mem_memoria: RAM_mem;

signal s_derechos_acceso: std_logic;
signal s_estado: tipoestado;
signal s_pet: tp_contro_e;

signal s_AF: std_logic;
signal s_est: st_estado;
signal s_control: tp_contro_cam_cntl;

signal s_peticion: tp_peticion;

signal s_esperado: st_bloque_dat;

signal inicializacion: std_logic;
signal parar: std_logic;
signal finaltraza: std_logic:= '0';

shared variable final : boolean := false;
signal ciclo: integer:= 0;

file S, S_pro_cons: text;

constant fichero: string := "../../../RESULTADOS/resultados_ejecucion.txt";
constant fichero_pro_cons: string := "../../../RESULTADOS/productor_consumidor.txt";

begin

ensamblado: jerarquia port map(reloj => reloj, pcero => pcero, pet_proc => peticion, resp_cache => respuesta, cache_lista => pet_listo);

-- captura de senyales internas al disenyo
-- cache: campos etqiuetas, estado y datos
	s_mem_etiq <= << signal .prueba_ensamblado.ensamblado.cache_bloqueante.cach_L2.cache.camino_datos_cache.etiquetas.memoria_etiquetas.campo_etiquetas: tp_m_ET >>;
	s_mem_estado <= << signal .prueba_ensamblado.ensamblado.cache_bloqueante.cach_L2.cache.camino_datos_cache.estado.campo_estado: tp_m_EST >>;
	s_mem_datos <= << signal .prueba_ensamblado.ensamblado.cache_bloqueante.cach_L2.cache.camino_datos_cache.datos.memoria_datos.campo_datos: tp_m_DAT >>;
-- memoria
	s_mem_memoria <= << signal .prueba_ensamblado.ensamblado.memoria.memoria_principal.memoria.memoria: RAM_mem >>;
-- controlador de cache: derechos de acceso, estado y peticion que se procesa
	s_derechos_acceso <= << signal .prueba_ensamblado.ensamblado.cache_bloqueante.cach_L2.cache.controlador_cache.derechos_acceso: std_logic >>;
	s_estado <= << signal .prueba_ensamblado.ensamblado.cache_bloqueante.cach_L2.cache.controlador_cache.estado: tipoestado >>;
--	s_pet <= << signal .prueba_ensamblado.ensa_ca_mem.cache.cach.cache_sin.contro.pet: tp_contro_e >>;
-- controlador de cache: senyales de entrada acierto/fallo, estado del bloque accedido
	s_AF <= << signal .prueba_ensamblado.ensamblado.cache_bloqueante.cach_L2.cache.camino_datos_cache.etiquetas.AF: std_logic >>;
	s_est <= << signal .prueba_ensamblado.ensamblado.cache_bloqueante.cach_L2.cache.camino_datos_cache.estado.DL: st_estado >>;
-- controlador de cache: senyales de control
	s_control <= << signal .prueba_ensamblado.ensamblado.cache_bloqueante.cach_L2.cache.controlador_cache.s_control: tp_contro_cam_cntl >>;
-- cache: peticion que procesa la cache
	s_peticion <= << signal .prueba_ensamblado.ensamblado.cache_bloqueante.cach_L2.cache.peticion: tp_peticion >>;


productor: process 
variable v_DIR: natural range 0 to tam_EspacioLogico;
variable v_DATO: natural range 0 to tam_palabra;
variable v_exp: std_logic; -- Identifica si la peticion que se envia es Pt o PtXl
begin
-- fichero resumen
 	file_open(S_pro_cons,fichero_pro_cons,write_mode); 
	cabecera_resumen (fichero_pro_cons);
	file_close(S_pro_cons);

-- fichero de traza     
	if (imprimir_traza = 1) then
		file_open(S,fichero,write_mode); 
		--cabecera_traza (fichero);
		file_close(S);
	end if;

-- puesta a cero
	proc_puesta_cero (reloj, pcero, peticion, pet_listo, ciclo, fichero_pro_cons);
	v_exp := '0';

-- inicio de peticiones
   -- Prueba con la peticion de inicio. Deja el contenedor en M tanto en L1 como en L2
   v_DIR := 0; 
	v_DATO := 3;
	inicio (reloj, peticion, pet_listo, v_DIR, v_DATO, ciclo, fichero_pro_cons);
	
	-- Llega una peticion PtX. Es acierto. Cambio de M a MNP
	Pescritura (reloj, peticion, pet_listo, v_DIR, v_DATO, ciclo, fichero_pro_cons);
	
	-- Llega una peticion Pt. Es a la direccion 0. L2 ha de suministrar el bloque. Cambio de estado de MNP a M
	Plectura (reloj, peticion, pet_listo, respuesta, s_esperado, v_DIR, v_DATO, ciclo, fichero_pro_cons, v_exp);
	
	-- Llega una peticion Pt. L2 no tiene el bloque por tanto emite una peticion Ptm a memoria y suministra el bloque a la L1. Estado L
	v_DIR := 6;
   Plectura (reloj, peticion, pet_listo, respuesta, s_esperado, v_DIR, v_DATO, ciclo, fichero_pro_cons, v_exp);
	
	-- Llega una peticion PtXl. Es acierto. Cambio de L a LNP
	v_exp := '1';
   Plectura (reloj, peticion, pet_listo, respuesta, s_esperado, v_DIR, v_DATO, ciclo, fichero_pro_cons, v_exp);
	
	-- De nuevo, peticion Pt a la @6. Es acierto en L2 y se suministra el dato. Cambio de LNP a L
	v_DIR := 6;
	v_exp := '0';
   Plectura (reloj, peticion, pet_listo, respuesta, s_esperado, v_DIR, v_DATO, ciclo, fichero_pro_cons, v_exp);
	
	-- Llega una peticion PtXl. Es acierto. Cambio de L a LNP
	v_exp := '1';
   Plectura (reloj, peticion, pet_listo, respuesta, s_esperado, v_DIR, v_DATO, ciclo, fichero_pro_cons, v_exp);
	
	-- Llega una peticion Pt. Reemplaza el bloque de la peticion anterior. Como se encuentra en LNP, no requiere actualizar memoria
	v_DIR := 38;
	v_exp := '0';
   Plectura (reloj, peticion, pet_listo, respuesta, s_esperado, v_DIR, v_DATO, ciclo, fichero_pro_cons, v_exp);
	
	-- Llega una peticion PtX a la direccion 0. Es acierto. Cambio de M a MNP
	v_DIR := 0;
	v_DATO := 3;
	Pescritura (reloj, peticion, pet_listo, v_DIR, v_DATO, ciclo, fichero_pro_cons);
	
	-- Peticion Pt a la @32, provocando el reemplazo del bloque almacenado en el contenedor 0. Esta en estado MNP. Ha de actualizarse memoria
	v_DIR := 32;
   v_exp := '0';
	Plectura (reloj, peticion, pet_listo, respuesta, s_esperado, v_DIR, v_DATO, ciclo, fichero_pro_cons, v_exp);

	no_hay_peticion (reloj, peticion, pet_listo, ciclo, fichero_pro_cons);
	no_hay_peticion (reloj, peticion, pet_listo, ciclo, fichero_pro_cons);

	interface_productor(reloj, pet_listo);

	report "prueba finalizada";

	parar <= '1';
	wait;       
end process;


consumidor: process is
variable v_s_peticion: tp_peticion;
variable esperado, consumo: st_bloque_dat;
variable ciclod:integer;
file S_pro_cons: text;
variable Lo, l : line;
begin
--	capturar valor esperado en una instruccion load (s_esperado)
	interface_productor(reloj, pet_listo);
	if peticion.acc = '1' and peticion.pe = '0' and peticion.ini = '0' then
		esperado := s_esperado; --ver

		interface_consumidor(reloj, respuesta.valido);

		consumo := respuesta.dato_leido;

-- Actualizar fichero. Instante en el cual se consume el valor del load 
		ciclod:= ciclo'delayed(0 fs);
		write(l, ciclod, right, 5);
		write (l, string'("consumo. valor"), right, 20+7); 
		hwrite(l, consumo, right, 6);
		write (l, string'("load  "), right, 8); 
		hwrite(l, s_peticion.dir, right, 6);
		file_open(S_pro_cons,fichero_pro_cons,append_mode); 
		writeline (S_pro_cons, l);
		file_close(S_pro_cons);

		if comprobar_load = 1 then
-- comprobacion del valor leido con el esperado
			if (respuesta.dato_leido /= esperado) then 
				assert false report "valor no esperado" severity warning;
				write(Lo, string'(", leido:   "));
				write(Lo, respuesta.dato_leido);
				write(Lo, string'(", esperado:   "));
				write(Lo, esperado);
				writeline(output, Lo);

				write(l, string'("valor no esperado "));
				write(l, string'(", leido:   "));
				write(l, respuesta.dato_leido);
				write(l, string'(", esperado:   "));
				write(l, esperado);
				file_open(S_pro_cons,fichero_pro_cons,append_mode); 
				writeline (S_pro_cons, l);
				file_close(S_pro_cons);
			end if;
		end if;
	end if;
end process;


--traza: if imprimir_traza = 1 generate
--impri_accesos: process
--
--variable v_peticion: tp_peticion;
--variable v_respuesta: tp_respuesta;
--variable v_pet_listo: st_cache_listo;
--
--variable v_derechos_acceso: std_logic;
--variable v_estado: tipoestado;
--variable v_pet: tp_contro_e;
--
--variable v_AF: std_logic;
--variable v_est: std_logic;
--variable v_control, v_control_actuacion: tp_contro_cam_cntl;
--
--variable v_s_peticion: tp_peticion;
--
--variable ciclod:integer;
--variable cnt, cnt_sigue: integer := 0;
--
--begin
--	wait until rising_edge(reloj);
--	v_pet_listo:= pet_listo'delayed(0 fs);
--	if ciclo >= 5 and finaltraza = '0' then
---- valor de las senyales en el instante previo al flanco ascendente
--		v_peticion:= peticion'delayed(0 fs);
--		v_respuesta:= respuesta'delayed(0 fs);
--		v_estado:= s_estado'delayed(0 fs);
--		v_pet:= s_pet'delayed(0 fs);
--		v_AF:= s_AF'delayed(0 fs);
--
--		v_est:= s_est'delayed(0 fs);
--
--		v_control:= s_control'delayed(0 fs);
--		v_s_peticion := s_peticion'delayed(0 fs);
--
--		ciclod:= ciclo'delayed(0 fs);
--
---- como los campos de cache y memoria no se actualizan en cada ciclo no es necesario "delayed"
--		impri_traza (v_pet_listo, v_s_peticion, v_peticion, v_AF, v_est, v_estado,
--					s_mem_etiq, s_mem_estado, s_mem_datos, s_mem_memoria,
--					v_control_actuacion,
-- 					ciclod, cnt, cnt_sigue, fichero);
--		v_control_actuacion := v_control;
--	end if;
--
--	if parar = '1' then
--		finaltraza <= '1';
--	end if;
--
--end process;
--end generate traza;


finalizar: process is
begin
	wait until parar = '1';
	final := true;
	if imprimir_cache = 1 then
		impri_cache(s_mem_etiq, s_mem_estado, s_mem_datos, fichero_pro_cons);
	end if;
	if imprimir_memoria = 1 then
		impri_memoria(s_mem_memoria, fichero_pro_cons);
	end if;
end process;


relojciclo: process  is
begin
  if final = false then
	reloj <= '0';
	wait for 40 ns;
	ciclo <= ciclo +1;
	reloj <= '1';
	wait for 40 ns;
	if pasoapaso = 1 then
		stop(0);
	end if;
  else
	wait;
  end if;
end process relojciclo;

end;
